* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 D RN SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vccd1 vssd1
XFILLER_54_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__050__A3 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_045_ net5 _003_ _018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_028_ net12 net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__044__A1 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output12_I net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_044_ net4 _016_ _017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_19_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_027_ net10 _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I io_in[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_043_ _010_ _002_ _016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__053__B net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_042_ _011_ _012_ _014_ _015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__038__A1 _008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput12 net12 io_out[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__029__A1 net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_041_ net2 _013_ _014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput13 net13 io_out[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__029__A2 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input1_I io_in[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_040_ _008_ _009_ _013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__038__A3 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__029__A3 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__037__I net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__040__A1 _008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__031__A1 net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__031__A2 net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__052__A1 net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I io_in[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__034__A1 net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 io_in[10] net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput2 io_in[11] net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput3 io_in[12] net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__055__A1 _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__056__RN _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__055__A2 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_056_ mod.flipflop1.d _000_ _001_ net8 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_7_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_039_ _008_ _009_ _010_ _002_ _012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 io_in[14] net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_80 io_oeb[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_51_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_055_ _000_ net9 _001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_038_ _008_ _009_ net2 _010_ _011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_70 io_oeb[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput6 io_in[15] net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_81 io_oeb[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_054_ _005_ _020_ _024_ _026_ mod.flipflop1.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_11_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_037_ net3 _010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I io_in[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_60 io_oeb[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_71 io_oeb[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput7 io_in[16] net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_82 io_oeb[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_053_ _005_ _025_ net12 _026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput10 io_in[19] net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_036_ net11 _009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 io_in[17] net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_50 io_oeb[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_72 io_oeb[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_61 io_oeb[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_83 io_oeb[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_052_ net7 _004_ _025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput11 io_in[9] net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_035_ net1 _008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__030__A1 net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__035__I net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_51 io_oeb[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_73 io_oeb[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_84 io_oeb[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput9 io_in[18] net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_40 io_out[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_62 io_oeb[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_051_ _005_ _021_ _022_ _023_ _024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_034_ net6 _006_ _007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__030__A2 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I io_in[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I io_in[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_41 io_out[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_85 io_oeb[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_30 io_out[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_52 io_oeb[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_63 io_oeb[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_74 io_oeb[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_050_ _008_ _009_ net2 _010_ _023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_033_ net5 _003_ _006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_31 io_out[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_20 io_out[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_86 io_oeb[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_42 io_out[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_53 io_oeb[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_75 io_oeb[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_64 io_oeb[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__033__A1 net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_032_ net7 _004_ _005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_65 io_oeb[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_54 io_oeb[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_32 io_out[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_21 io_out[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_43 io_out[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_76 io_oeb[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_87 io_oeb[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_031_ net6 net5 _003_ _004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_3_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_22 io_out[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_77 io_oeb[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_33 io_out[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_44 io_out[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_55 io_oeb[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_66 io_oeb[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_030_ net3 net4 _002_ _003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_3_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_34 io_out[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_56 io_oeb[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_45 io_out[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_23 io_out[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_67 io_oeb[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_78 io_oeb[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__045__A1 net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_68 io_oeb[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_35 io_out[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_79 io_oeb[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_46 io_out[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_24 io_out[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_57 io_oeb[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_36 io_out[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_25 io_out[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_47 io_out[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_14 io_out[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_69 io_oeb[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_58 io_oeb[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input9_I io_in[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_59 io_oeb[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_37 io_out[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_48 io_out[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_15 io_out[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_26 io_out[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__039__A1 _008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_38 io_out[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_49 io_out[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_16 io_out[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_27 io_out[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_17 io_out[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_39 io_out[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_28 io_out[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input7_I io_in[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_18 io_out[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_29 io_out[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__028__I net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_049_ _017_ _018_ _015_ _022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_19 io_out[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__036__I net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_048_ _017_ _018_ _015_ _021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_19_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__056__CLK net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__050__A1 _008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__041__A1 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__032__A1 net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_047_ _007_ _015_ _019_ _020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_34_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input5_I io_in[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_046_ _017_ _018_ _019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_029_ net1 net11 net2 _002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

